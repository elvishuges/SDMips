
`timescale 1ns/10ps

module somador_pc_tb;


reg [31:0] op_1;
wire [31:0] resul_soma;


somador_pc dut(.op_1(op_1),.resul_soma(resul_soma));

initial
begin



op_1 = 32'b00000000000000000000000000000000;
#0.1;
op_1 = 32'b00000000000000000000000000000001;
#0.1;
op_1 = 32'b00000000000000000000000000000010;
#0.1;
op_1 = 32'b00000000000000000000000000000011;
#0.1;
op_1 = 32'b00000000000000000000000000000100;


end

endmodule
